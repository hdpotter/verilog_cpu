module if_id(
    input logic [31:0] instr_in,
    output logic [31:0] instr_out,

    input clk,
    input rst
);

always @(posedge clk) begin
    if(!rst) begin
        instr_out <= instr_in;
    end else begin
        instr_out <= 32'h00000013; //nop on reset
    end
end

endmodule